library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


use IEEE.NUMERIC_STD.ALL;


entity ROM is
  Port (
         A: in std_logic_vector(9 downto 0);
         D: out std_logic_vector(15 downto 0);
         en_ROM:in std_logic ;
			clk:in std_logic);
end ROM;

architecture Behavioral of ROM is

    
    type rom_type is array(0 to 63) of std_logic_vector(15 downto 0);
    
    constant program: rom_type:=(
		  "0001100000000000",
		  "0000010000000000",
		  "0001010000000000",
		  "0001010000000000",
		  "0001010000000000",
		  "0001010000000000",
		  "0001010000000000",
		  "1000000000000000",
		  "0010000000000000",
		  "0010010000000000",
		  "0010010000000000",
		  "0011100000000000",
		  "0011100000000000",
		  "0011100000000000",
		  "0011110000000000",
		  "0011110000000000",
		  "0011110000000000",
		  "0001100000000000",
		  "0010000000000000",
		  "0010000000000000",
		  "0010000000000000",
		  "0010000000000000",
		  "0010000000000000", 
		  "0010000000000000",
		  "0010000000000000",
        "0010000000000000",
        "0010000000000000",
        "0010010000000000",
        "0010010000000000",
        "0010010000000000",
        "0010010000000000",
        "0010010000000000",
        "0010010000000000",
        "0010000000000000",
        "0010000000000000",
        "0010000000000000",
        "0010000000000000",
        "0010000000000000",
        "0010000000000000",
        "0010000000000000",
        "0010000000000000",
        "0010000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000"
    );
begin
		process(clk)
		begin
				if(rising_edge(clk) and en_rom = '1') then		
					D<=program(to_integer(unsigned(A)));
			   end if;
		end process;
end Behavioral;